LAB1

.LIB "EVAL.LIB"

V1 1 0 DC 1
D1 1 0 D1N4148

.DC V1 0 1 0.01
.TEMP 0 25 50
.PROBE
.END