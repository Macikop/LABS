Kolos1

R1 4 3 30
R2 4 5 6
R3 2 7 8
R4 4 0 30
R5 6 4 15
R6 2 1 40

L1 1 0 10u
C1 6 0 1u

V1 2 3 30
V2 0 5 200
V3 0 7 60

VA 2 6 0

H1 4 0 VA 20

.DC V1 30 30 1
.TF V(2) V1
.PRINT DC W(V1) W(V2) W(V3) I(R6) W(R6) V(2)
.END