Lab4

R1 3 0 5
R2 1 0 5

L1 5 2 0.159
C1 4 2 1.59M

V1 2 3 AC 20
V2 1 4 AC 10 -90
V3 1 5 AC 10 90
I1 0 1 AC 5

.AC LIN 1 10 10
.PRINT AC VR(L1) VI(L1) VR(C1) VI(C1) VM(2,3) VP(2,3)
.END
Lab4

R1 3 0 5
R2 1 0 5

L1 5 6 0.159
RL 2 6 1N
C1 4 2 1.59M

V1 2 3 AC 20
V2 1 4 AC 10 -90
V3 1 5 AC 10 90
I1 0 1 AC 5

VX 2 4 0

.AC LIN 1 10 10
.PRINT AC IM(VX) IP(VX)
.END