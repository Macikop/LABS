Lab7

.MODEL VSW VSWITCH RON=1m ROFF=1G VOFF=0 VON=1

VT 4 0 PULSE(0 1 1m)
RT 4 0 10

C1 1 0 1u IC=5
R1 2 1 20
S1 3 2 4 0 VSW
L1 3 0 10m

.TRAN 0 10m 0 100n
.PROBE
.END