KOLOS A

.LIB "EVAL_TOS.LIB"

.PARAM CURRENT = 1U
.PARAM AMP = 1.17M
.PARAM W = 48.7U
VP VDD 0 DC 5

*VIN IN 0 DC 707.034M AC 1 SIN(707.034M, {AMP}, 100K)
VIN IN 0 PULSE(0 5 10N)
IREF GATES 0 {CURRENT}

M1 1 GATES VDD VDD PMOS0P5 W=15U L=0.3U
M2 2 GATES VDD VDD PMOS0P5 W=15U L=0.3U
M3 GATES GATES 1 VDD PMOS0P5 W=15U L=0.3U
M4 OUT GATES 2 VDD PMOS0P5 W=15U L=0.3U

M5 OUT IN 0 0 NMOS0P5 W={W} L=0.3U

C1 OUT 0 200P
*.DC VIN 0 1 100u
*.STEP LIN PARAM CURRENT 0.1U 100U 0.1U
*.DC VIN 700M 710M 100N
*.AC DEC 10 1 1GHZ 
*.TRAN 0 100U 0 100N
*.STEP LIN PARAM AMP 100U 10M 10U
*.FOUR 100K V[OUT]
*.TF V[OUT] VIN

.TRAN 0 50N 0 1N
*.STEP LIN PARAM W 30U 60U 0.1U
.PROBE
.END

;iref = 0.1u kv = -7k
