Lab4

V1 1 0 SIN(1 1 1kHz)

R1 1 2 1k
C1 2 0 159n

.TRAN 0 10m 0 10n
.FOUR 1kHz V(2)
.PROBE
.END