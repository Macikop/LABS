KOLOS2A

.LIB "EVAL_TOS.LIB"

.PARAM CAP = 520U

V1 VX 0 SIN(0 169.2 60)

RX VX VIN 1P

XTRAFO VIN 0 OUTP 0 OUTN TX_I

D1 OUTP 1 D1N4148
D2 OUTN 1 D1N4148

C1 1 0 {CAP}
R1 1 2 191
*XZENER 0 2 ZENER_I

RL 2 0 150

.TRAN 0 5 4.0 1M
.STEP LIN PARAM CAP 20M 20M 1M
.PROBE
.END
