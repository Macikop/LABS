KOLOS2

.LIB "EVAL_TOS.LIB"

.PARAM CAP = 500U

V1 9 0 SIN(0 84.85 60)
RV 9 1 1N

XTRAFO 1 0 2 3 TX_II

D1 2 4 D1N4148
D2 0 3 D1N4148
D3 3 4 D1N4148
D4 0 2 D1N4148

C1 4 0 {CAP}
R1 4 5 200
XZ 0 5 ZENER_II
RL 5 0 1K

.STEP LIN PARAM CAP 1M 50M 1M

.TRAN 0 10 9 1M
.PROBE

.END