LAB5

.LIB "EVAL.LIB"

.MODEL INZ1 D IS=100 N=0.01
.MODEL INZ2 D IS=100 N=1.679

.SUBCKT ZENER ANODE CATODE

	RZ ANODE 1 20
	VZ 2 1 6.7
	D1 CATODE 2 INZ1
	D2 ANODE CATODE INZ2

.ENDS


V1 1 0 10
R1 1 2 1k
XZ 0 2 ZENER
RL 2 0 2K

.DC LIN V1 9 11 0.1
.PROBE
.END 