Lab1

.LIB "EVAL.LIB"

VCC VCC 0 15
VEE 0 VEE 15

V_P IN_P 0 0 AC 1
V_N IN_N 0 0

XOPAMP IN_P IN_N VCC VEE OUT UA741

.DC V_P -0.01 0.01 0.0001
.AC DEC 10 1HZ 10MEGHZ

.TF V[OUT] V_P

.PROBE
.END