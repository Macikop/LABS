Lab1

V1 1 0 AC 1

R1 1 2 1k
C1 2 0 159n

.AC DEC 100 1 1MEG

.PROBE
.END