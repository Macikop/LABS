Lab5

R1 2 1 10

L1 3 6 3.183M
RL 5 6 1P

C1 3 4 31.83U

VX 4 1 0

V1 2 0 AC 20 90
V2 1 0 AC 5 0
V3 5 0 AC 20

F1 2 1 VX 2
E1 1 3 2 1 3

.AC LIN 1 500 500 
.PRINT AC IM(V1) IM(V2) IM(V3) IP(V1) IP(V2) IP(V3)
.END