LAB4

.LIB "EVAL.LIB"

.PARAM AMP = 0

VIN 1 0 AC {AMP}
R1 1 2 1K

D1 2 3 D1N4148
V1 3 0 DC 5

D2 4 2 D1N4148
V2 0 4 DC 4

*.STEP LIN PARAM AMP -8 8 1

.DC VIN -20 20 1

.PROBE

.END