KOLOS B

.LIB "EVAL_TOS.LIB"

.PARAM RES = 100K
.PARAM AMP = 5.8M
.PARAM W = 100U

VP VDD 0 DC 5

M1 1 1 VDD VDD PMOS0P5 W=10U L=0.5U
M2 OUT 1 VDD VDD PMOS0P5 W=10U L=0.5U

M3 2 2 0 0 NMOS0P5 W=10U L=0.5U
M4 OUT IN 0 0 NMOS0P5 W={W} L=0.5U

R1 1 2 {RES}

*VIN IN 0 DC 736.012M AC 1 SIN(736.012M, {AMP}, 100K)
VIN IN 0 PULSE(5 0 1U)
C1 OUT 0 2N
*KV=-260.472
*.DC VIN 0 5 100U
*.STEP LIN PARAM RES 1K 100K 1K

*.DC VIN 700M 750M 1U
*.AC DEC 10 1 1G
.TRAN 0 20U 0 1N
*.STEP LIN PARAM AMP 100U 10M 100U
*.FOUR 100K V[OUT]

.STEP LIN PARAM W 50U 150U 1U

.PROBE
.END