Lab3

R1 4 0 39
R2 5 0 18
R3 2 1 72

Vx 3 5 0

V1 4 3 10
I1 0 1 1.6

H1 3 2  Vx 40

.DC V1 10 10 1

.PRINT DC V(H1) I(H1) W(H1) V(R2) I(R2) W(R2) V(0,2)
.TF V(0,2) V1
.END