Lab2

.PARAM RESISTANCE = 100

V1 1 0 AC 1

R1 1 2 {RESISTANCE}
C1 2 0 159n

.AC DEC 2 1 100K
.STEP DEC PARAM RESISTANCE 100 10K 2 
.PROBE
.END