Lab3

.MODEL RT RES R=1 TC1=0.01
.MODEL CT CAP C=1 TC1=-0.002

V1 1 0 AC 1

R1 1 2 RT 1k
C1 2 0 CT 159n

.AC DEC 10 1 1MEG
.TEMP 0 40 80 120
.PROBE
.END