LAB3

.LIB "EVAL.LIB"

.PARAM OFFSET = 0

V1 1 0 SIN({OFFSET} 10 1) 
D1 1 2 D1N4148
R1 2 0 1K
c1 2 0 39m

.STEP LIN PARAM OFFSET 9 10 0.1
.TRAN 0 2 0 1M
.FOUR 1 V(2)
.PROBE

.END