Lab6

V1 9 0 AC 200
RTR 9 1 1P

L1 1 0 0.239
L2 2 0 0.159
KTR L1 L2 1

R1 3 2 0.333
C1 4 3 0.477

L3 4 0 0.08
R2 4 0 1

R3 5 4 1
L4 6 5 0.159
C2 6 0 0.08

.AC DEC 100 0.1 10
.PROBE
.END
 