Lab2

.LIB "EVAL.LIB"

V_P IN_P 0 PULSE(0 10)

VCC VCC 0 15
VEE 0 VEE 15

XOPAMP IN_P OUT VCC VEE OUT UA741

R1 OUT 0 2K
C1 OUT 0 100P

.TRAN 0 30U 0 10N

.PROBE
.END