KOLOS C

.LIB "EVAL_TOS.LIB"

VIN IN 0 DC 3
VP VDD 0 DC 5

M1 VDD IN 0 0 PMOS0P5

.DC VP 0 5 0.1
.PROBE
.END