Lab8

.MODEL VSW VSWITCH RON=1m ROFF=1G VOFF=0 VON=1
.MODEL VSWn VSWITCH RON=1m ROFF=1G VOFF=1 VON=0

VT 6 0 PULSE(0 1 0.5m)
RT 6 0 10

C1 1 0 100n
R1 2 1 10
S1 2 4 6 0 VSW
L1 4 0 1m
S2 3 4 6 0 VSWn
R2 5 3 2k
V1 5 0 2

.TRAN 0 2m 0 10n
.PROBE
.END