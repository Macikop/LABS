Lab1

R1 1 2 80
R2 3 1 70
R3 2 0 60
R4 3 0 90

V1 2 3 2
I1 0 1 0.2

.DC V1 2 2 1
.OP
.PRINT DC V(R3) I(R4)
.END