Lab2

R1 2 1 100
R2 3 2 40
R3 0 3 170
R4 1 3 70
R5 2 0 50
R6 1 0 20

I1 0 1 1

.TF V(1) I1

.END