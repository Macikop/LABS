LAB2

.LIB "EVAL.LIB"

V1 1 0 DC 10 AC 0.1 
R1 1 2 1K
D1 2 0 D1N4148



.SENS V(2)
.AC LIN 1 1KHZ 1KHZ
.PRINT AC V(2) I(D1)
.END